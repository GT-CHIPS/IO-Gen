* Momentum eesofbbs_64 12.00 (*) built: Jan 14 2016
**************************************************
*.LIB Case1_5mm

*bbspice subcircuit with consecutive port numbers.

.SUBCKT bbspice_subckt	  port_1  port_2  port_3  port_4  port_5  port_6  gnd_0

* PORT_1
vi_1	port_1	_net_1	0.00000000000000e+000
vb_1	_net_4	_net_5	0.00000000000000e+000
R_Z0_1 	_net_1 	_net_2 	5.00000000000000e+001	NOISE=0
H_b_1	_net_2	gnd_0	vb_1	1.41421356237310e+001
E_v_1	_net_3	gnd_0	port_1	gnd_0	7.07106781186548e-002
H_i_1	_net_4	_net_3	vi_1	3.53553390593274e+000


G_POLE_port1_port1_p1 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	4.82651001152243e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port1_port1_p2 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	1.43365773872699e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port1_port1_p3 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	1.27519591890766e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port1_port1_p4 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	1.78504427429108e+010 	1.09642668997895e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port1_port2_p1 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	5.07966415829811e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port1_port2_p2 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	1.36216706913382e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port1_port2_p3 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	-4.60790790353513e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port1_port2_p4 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	4.38884155596893e+010 	6.89451147614233e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port1_port3_p1 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.80216185006337e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port1_port3_p2 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	5.35189742199792e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port1_port3_p3 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	4.00206027869048e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port1_port3_p4 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	7.73070058654280e+010 	-1.17024417578864e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port1_port4_p1 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.58633040522622e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port1_port4_p2 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	4.84953165965305e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port1_port4_p3 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	4.29888109132133e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port1_port4_p4 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	-3.70033906165474e+010 	3.94149523980163e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port1_port5_p1 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	1.23276077058375e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port1_port5_p2 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	-8.87859999207361e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port1_port5_p3 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	5.98967119572984e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port1_port5_p4 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	-8.54319029331276e+009 	1.57270206364419e+012 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port1_port6_p1 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	1.30161532017439e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port1_port6_p2 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.36551308651680e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port1_port6_p3 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	2.25579848301703e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port1_port6_p4 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-2.32724553023585e+010 	-3.48274187899991e+009 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010

* PORT_2
vi_2	port_2	_net_6	0.00000000000000e+000
vb_2	_net_9	_net_10	0.00000000000000e+000
R_Z0_2 	_net_6 	_net_7 	5.00000000000000e+001	NOISE=0
H_b_2	_net_7	gnd_0	vb_2	1.41421356237310e+001
E_v_2	_net_8	gnd_0	port_2	gnd_0	7.07106781186548e-002
H_i_2	_net_9	_net_8	vi_2	3.53553390593274e+000


G_POLE_port2_port1_p1 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	5.07966415829811e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port2_port1_p2 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	1.36216706913382e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port2_port1_p3 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	-4.60790790353513e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port2_port1_p4 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	4.38884155596893e+010 	6.89451147614233e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port2_port2_p1 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	4.70171024140511e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port2_port2_p2 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	1.35178766112809e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port2_port2_p3 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	1.71259831242169e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port2_port2_p4 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	1.53569391409913e+010 	9.45130118488432e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port2_port3_p1 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.62894598098968e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port2_port3_p2 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	5.25669383770125e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port2_port3_p3 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	3.96014568586686e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port2_port3_p4 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	-3.42835156227121e+010 	3.98697616700504e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port2_port4_p1 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.59463428021032e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port2_port4_p2 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	5.43083138709749e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port2_port4_p3 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	3.72263180693263e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port2_port4_p4 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	7.86838289904377e+010 	-1.08926430533806e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port2_port5_p1 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	1.25558482067280e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port2_port5_p2 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.33022191200120e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port2_port5_p3 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	1.99594471815688e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port2_port5_p4 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-2.11892074953218e+010 	-3.64528604766552e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port2_port6_p1 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	1.11054515107879e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port2_port6_p2 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	-8.00868530033351e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port2_port6_p3 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	5.94147438011760e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port2_port6_p4 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	-8.95172625554374e+009 	1.54609473603977e+012 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010

* PORT_3
vi_3	port_3	_net_11	0.00000000000000e+000
vb_3	_net_14	_net_15	0.00000000000000e+000
R_Z0_3 	_net_11 	_net_12 	5.00000000000000e+001	NOISE=0
H_b_3	_net_12	gnd_0	vb_3	1.41421356237310e+001
E_v_3	_net_13	gnd_0	port_3	gnd_0	7.07106781186548e-002
H_i_3	_net_14	_net_13	vi_3	3.53553390593274e+000


G_POLE_port3_port1_p1 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-3.80216185006337e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port3_port1_p2 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	5.35189742199792e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port3_port1_p3 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	4.00206027869048e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port3_port1_p4 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	7.73070058654280e+010 	-1.17024417578864e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port3_port2_p1 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	-3.62894598098968e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port3_port2_p2 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	5.25669383770125e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port3_port2_p3 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	3.96014568586686e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port3_port2_p4 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	-3.42835156227121e+010 	3.98697616700504e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port3_port3_p1 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	3.75199167477779e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port3_port3_p2 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	1.73612135115996e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port3_port3_p3 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	1.97526129147995e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port3_port3_p4 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	3.05498768198560e+010 	-4.22057859723639e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port3_port4_p1 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	3.90647400886121e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port3_port4_p2 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	1.69033626026053e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port3_port4_p3 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.37063715687125e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port3_port4_p4 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	3.01731483809985e+010 	-6.37369292218294e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port3_port5_p1 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-3.66965707626241e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port3_port5_p2 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	4.72792781332274e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port3_port5_p3 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	4.28473533220259e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port3_port5_p4 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	7.45897157746694e+010 	-1.30679924449104e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port3_port6_p1 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	-3.51166077095456e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port3_port6_p2 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	4.59743892618759e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port3_port6_p3 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	4.37887503333026e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port3_port6_p4 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	-3.71385747226743e+010 	3.98280790737238e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010

* PORT_4
vi_4	port_4	_net_16	0.00000000000000e+000
vb_4	_net_19	_net_20	0.00000000000000e+000
R_Z0_4 	_net_16 	_net_17 	5.00000000000000e+001	NOISE=0
H_b_4	_net_17	gnd_0	vb_4	1.41421356237310e+001
E_v_4	_net_18	gnd_0	port_4	gnd_0	7.07106781186548e-002
H_i_4	_net_19	_net_18	vi_4	3.53553390593274e+000


G_POLE_port4_port1_p1 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	-3.58633040522622e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port4_port1_p2 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	4.84953165965305e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port4_port1_p3 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	4.29888109132133e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port4_port1_p4 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	-3.70033906165474e+010 	3.94149523980163e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port4_port2_p1 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-3.59463428021032e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port4_port2_p2 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	5.43083138709749e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port4_port2_p3 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	3.72263180693263e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port4_port2_p4 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	7.86838289904377e+010 	-1.08926430533806e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port4_port3_p1 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	3.90647400886121e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port4_port3_p2 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	1.69033626026053e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port4_port3_p3 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.37063715687125e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port4_port3_p4 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	3.01731483809985e+010 	-6.37369292218294e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port4_port4_p1 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	3.53154832834560e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port4_port4_p2 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	1.67531610670302e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port4_port4_p3 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	1.84489093055063e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port4_port4_p4 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	3.78073847937061e+010 	6.64746038742487e+009 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port4_port5_p1 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	-3.49716223913043e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port4_port5_p2 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	4.33112593601920e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port4_port5_p3 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	4.68404515034247e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port4_port5_p4 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	-3.95108495144563e+010 	3.96438068993448e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port4_port6_p1 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-3.52488956553082e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port4_port6_p2 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	4.95624487238406e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port4_port6_p3 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	4.03077533860790e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port4_port6_p4 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	7.61738696743440e+010 	-1.23043267666664e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010

* PORT_5
vi_5	port_5	_net_21	0.00000000000000e+000
vb_5	_net_24	_net_25	0.00000000000000e+000
R_Z0_5 	_net_21 	_net_22 	5.00000000000000e+001	NOISE=0
H_b_5	_net_22	gnd_0	vb_5	1.41421356237310e+001
E_v_5	_net_23	gnd_0	port_5	gnd_0	7.07106781186548e-002
H_i_5	_net_24	_net_23	vi_5	3.53553390593274e+000


G_POLE_port5_port1_p1 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	1.23276077058375e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port5_port1_p2 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	-8.87859999207361e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port5_port1_p3 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	5.98967119572984e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port5_port1_p4 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	-8.54319029331276e+009 	1.57270206364419e+012 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port5_port2_p1 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	1.25558482067280e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port5_port2_p2 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.33022191200120e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port5_port2_p3 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	1.99594471815688e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port5_port2_p4 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.11892074953218e+010 	-3.64528604766552e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port5_port3_p1 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.66965707626241e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port5_port3_p2 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	4.72792781332274e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port5_port3_p3 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	4.28473533220259e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port5_port3_p4 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	7.45897157746694e+010 	-1.30679924449104e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port5_port4_p1 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.49716223913043e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port5_port4_p2 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	4.33112593601920e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port5_port4_p3 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	4.68404515034247e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port5_port4_p4 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	-3.95108495144563e+010 	3.96438068993448e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port5_port5_p1 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	4.71864334079048e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port5_port5_p2 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	1.45646764051475e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port5_port5_p3 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	1.15706620489494e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port5_port5_p4 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	1.04611179284158e+010 	2.29291929668141e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port5_port6_p1 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	4.95178360606320e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port5_port6_p2 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	1.41289075600869e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port5_port6_p3 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	-4.65097484256553e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port5_port6_p4 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	4.40262640237738e+010 	6.74341993270601e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010

* PORT_6
vi_6	port_6	_net_26	0.00000000000000e+000
vb_6	_net_29	_net_30	0.00000000000000e+000
R_Z0_6 	_net_26 	_net_27 	5.00000000000000e+001	NOISE=0
H_b_6	_net_27	gnd_0	vb_6	1.41421356237310e+001
E_v_6	_net_28	gnd_0	port_6	gnd_0	7.07106781186548e-002
H_i_6	_net_29	_net_28	vi_6	3.53553390593274e+000


G_POLE_port6_port1_p1 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	1.30161532017439e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port6_port1_p2 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.36551308651680e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port6_port1_p3 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	2.25579848301703e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port6_port1_p4 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.32724553023585e+010 	-3.48274187899991e+009 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port6_port2_p1 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	1.11054515107879e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port6_port2_p2 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	-8.00868530033351e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port6_port2_p3 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	5.94147438011760e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port6_port2_p4 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	-8.95172625554374e+009 	1.54609473603977e+012 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port6_port3_p1 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.51166077095456e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port6_port3_p2 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	4.59743892618759e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port6_port3_p3 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	4.37887503333026e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port6_port3_p4 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	-3.71385747226743e+010 	3.98280790737238e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port6_port4_p1 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.52488956553082e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port6_port4_p2 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	4.95624487238406e+009 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port6_port4_p3 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	4.03077533860790e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port6_port4_p4 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	7.61738696743440e+010 	-1.23043267666664e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port6_port5_p1 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	4.95178360606320e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port6_port5_p2 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	1.41289075600869e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port6_port5_p3 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	-4.65097484256553e+010 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port6_port5_p4 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	4.40262640237738e+010 	6.74341993270601e+010 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010
G_POLE_port6_port6_p1 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	4.53254019982106e+009 / 1.0 	1.91232730987567e+010 , 0.0
G_POLE_port6_port6_p2 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	1.45546830705480e+010 / 1.0 	4.30546876565498e+010 , 0.0
G_POLE_port6_port6_p3 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	9.25902133569766e+009 / 1.0 	1.16067082520069e+011 , 0.0
G_POLE_port6_port6_p4 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	2.03528539297943e+010 	1.79051716569122e+011 , 0.0 / 1.0 	1.92717631689730e+011 , -1.08212641732223e+010


.ENDS  bbspice_subckt
***************************************


***************************************
* S-based subckt

 
*bbspice subcircuit with external port numbers.

*.SUBCKT bbspice_Case1_5mm		1 	2 	3 	4 	5 	6 	0 
*
*x_ 	1 	2 	3 	4 	5 	6 	0 	bbspice_Case1_5mm_subckt
*
*.ENDS  bbspice_Case1_5mm
****************************************
*.ENDL
