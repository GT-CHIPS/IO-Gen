* Momentum eesofbbs_64 12.00 (*) built: Jan 14 2016
**************************************************
*.LIB Case2_1mm

*bbspice subcircuit with consecutive port numbers.

.SUBCKT bbspice_subckt	  port_1  port_2  port_3  port_4  port_5  port_6  gnd_0

* PORT_1
vi_1	port_1	_net_1	0.00000000000000e+000
vb_1	_net_4	_net_5	0.00000000000000e+000
R_Z0_1 	_net_1 	_net_2 	5.00000000000000e+001	NOISE=0
H_b_1	_net_2	gnd_0	vb_1	1.41421356237310e+001
E_v_1	_net_3	gnd_0	port_1	gnd_0	7.07106781186548e-002
H_i_1	_net_4	_net_3	vi_1	3.53553390593274e+000


G_POLE_port1_port1_p1 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-4.21356140029010e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port1_port1_p2 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.68216980956289e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port1_port1_p3 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.80329540308982e+010 	-2.97199404074539e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port1_port2_p1 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	3.77304505895140e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port1_port2_p2 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	2.91529389767688e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port1_port2_p3 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	-4.81726085027752e+010 	-8.42610274937035e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port1_port3_p1 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.01573900209750e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port1_port3_p2 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.84293401653714e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port1_port3_p3 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	9.59429887869213e+010 	3.18045127430416e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port1_port4_p1 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	2.19245915570141e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port1_port4_p2 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	1.34846695961521e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port1_port4_p3 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.74715039991097e+010 	1.49573845215966e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port1_port5_p1 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	5.71375830615799e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port1_port5_p2 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.12709850673771e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port1_port5_p3 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	5.34971913516873e+010 	3.85196714718207e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port1_port6_p1 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	-5.42018826291288e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port1_port6_p2 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	1.03434107472532e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port1_port6_p3 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-3.41448603628818e+009 	5.79437145226641e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010

* PORT_2
vi_2	port_2	_net_6	0.00000000000000e+000
vb_2	_net_9	_net_10	0.00000000000000e+000
R_Z0_2 	_net_6 	_net_7 	5.00000000000000e+001	NOISE=0
H_b_2	_net_7	gnd_0	vb_2	1.41421356237310e+001
E_v_2	_net_8	gnd_0	port_2	gnd_0	7.07106781186548e-002
H_i_2	_net_9	_net_8	vi_2	3.53553390593274e+000


G_POLE_port2_port1_p1 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	3.77304505895140e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port2_port1_p2 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	2.91529389767688e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port2_port1_p3 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	-4.81726085027752e+010 	-8.42610274937035e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port2_port2_p1 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-4.17872123276859e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port2_port2_p2 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.73968225556237e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port2_port2_p3 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.84498523898096e+010 	-2.93364090677653e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port2_port3_p1 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	2.19205036644677e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port2_port3_p2 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	1.35553600329468e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port2_port3_p3 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	-1.73952766219242e+010 	1.50600694815122e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port2_port4_p1 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.98594530974919e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port2_port4_p2 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.87581176625292e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port2_port4_p3 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	9.56701298865562e+010 	3.22018444370521e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port2_port5_p1 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	-5.39708544752101e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port2_port5_p2 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	1.03213272899589e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port2_port5_p3 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-3.43653656434887e+009 	5.75137884300703e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port2_port6_p1 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	5.80105329516571e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port2_port6_p2 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.13978752587401e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port2_port6_p3 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	5.33721279797821e+010 	3.88208408411310e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010

* PORT_3
vi_3	port_3	_net_11	0.00000000000000e+000
vb_3	_net_14	_net_15	0.00000000000000e+000
R_Z0_3 	_net_11 	_net_12 	5.00000000000000e+001	NOISE=0
H_b_3	_net_12	gnd_0	vb_3	1.41421356237310e+001
E_v_3	_net_13	gnd_0	port_3	gnd_0	7.07106781186548e-002
H_i_3	_net_14	_net_13	vi_3	3.53553390593274e+000


G_POLE_port3_port1_p1 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.01573900209750e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port3_port1_p2 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.84293401653714e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port3_port1_p3 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	9.59429887869213e+010 	3.18045127430416e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port3_port2_p1 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	2.19205036644677e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port3_port2_p2 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	1.35553600329468e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port3_port2_p3 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.73952766219242e+010 	1.50600694815122e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port3_port3_p1 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-4.88960410245129e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port3_port3_p2 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.67647001385408e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port3_port3_p3 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	4.03519597432032e+009 	1.53590623598872e+012 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port3_port4_p1 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	4.56212334493075e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port3_port4_p2 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	3.76609791889661e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port3_port4_p3 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	-3.29810049370898e+010 	-1.20910735378331e+012 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port3_port5_p1 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.99976607634523e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port3_port5_p2 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.84540716384569e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port3_port5_p3 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	9.61176083178391e+010 	3.17567816111629e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port3_port6_p1 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	2.16666961187778e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port3_port6_p2 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	1.38148736428337e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port3_port6_p3 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.75646416707469e+010 	1.50395977768986e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010

* PORT_4
vi_4	port_4	_net_16	0.00000000000000e+000
vb_4	_net_19	_net_20	0.00000000000000e+000
R_Z0_4 	_net_16 	_net_17 	5.00000000000000e+001	NOISE=0
H_b_4	_net_17	gnd_0	vb_4	1.41421356237310e+001
E_v_4	_net_18	gnd_0	port_4	gnd_0	7.07106781186548e-002
H_i_4	_net_19	_net_18	vi_4	3.53553390593274e+000


G_POLE_port4_port1_p1 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	2.19245915570141e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port4_port1_p2 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	1.34846695961521e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port4_port1_p3 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.74715039991097e+010 	1.49573845215966e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port4_port2_p1 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.98594530974919e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port4_port2_p2 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.87581176625292e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port4_port2_p3 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	9.56701298865562e+010 	3.22018444370521e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port4_port3_p1 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	4.56212334493075e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port4_port3_p2 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	3.76609791889661e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port4_port3_p3 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	-3.29810049370898e+010 	-1.20910735378331e+012 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port4_port4_p1 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-4.92824178675756e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port4_port4_p2 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.64678217427534e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port4_port4_p3 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	4.30537804275134e+009 	1.43403032398363e+012 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port4_port5_p1 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	2.16724146313207e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port4_port5_p2 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	1.37620130583179e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port4_port5_p3 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.76305730291661e+010 	1.49554659268587e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port4_port6_p1 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.96964053709550e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port4_port6_p2 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.88462510318307e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port4_port6_p3 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	9.57369477165946e+010 	3.22486483351622e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010

* PORT_5
vi_5	port_5	_net_21	0.00000000000000e+000
vb_5	_net_24	_net_25	0.00000000000000e+000
R_Z0_5 	_net_21 	_net_22 	5.00000000000000e+001	NOISE=0
H_b_5	_net_22	gnd_0	vb_5	1.41421356237310e+001
E_v_5	_net_23	gnd_0	port_5	gnd_0	7.07106781186548e-002
H_i_5	_net_24	_net_23	vi_5	3.53553390593274e+000


G_POLE_port5_port1_p1 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	5.71375830615799e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port5_port1_p2 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.12709850673771e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port5_port1_p3 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	5.34971913516873e+010 	3.85196714718207e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port5_port2_p1 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	-5.39708544752101e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port5_port2_p2 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	1.03213272899589e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port5_port2_p3 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-3.43653656434887e+009 	5.75137884300703e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port5_port3_p1 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.99976607634523e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port5_port3_p2 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.84540716384569e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port5_port3_p3 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	9.61176083178391e+010 	3.17567816111629e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port5_port4_p1 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	2.16724146313207e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port5_port4_p2 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	1.37620130583179e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port5_port4_p3 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.76305730291661e+010 	1.49554659268587e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port5_port5_p1 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-4.14345576733323e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port5_port5_p2 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.75605301342350e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port5_port5_p3 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.65022603146141e+010 	-3.28624712878193e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port5_port6_p1 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	3.74108139465422e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port5_port6_p2 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	2.92153191949078e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port5_port6_p3 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	-4.74723615989712e+010 	-8.54982158167148e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010

* PORT_6
vi_6	port_6	_net_26	0.00000000000000e+000
vb_6	_net_29	_net_30	0.00000000000000e+000
R_Z0_6 	_net_26 	_net_27 	5.00000000000000e+001	NOISE=0
H_b_6	_net_27	gnd_0	vb_6	1.41421356237310e+001
E_v_6	_net_28	gnd_0	port_6	gnd_0	7.07106781186548e-002
H_i_6	_net_29	_net_28	vi_6	3.53553390593274e+000


G_POLE_port6_port1_p1 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	-5.42018826291288e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port6_port1_p2 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	1.03434107472532e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port6_port1_p3 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-3.41448603628818e+009 	5.79437145226641e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port6_port2_p1 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	5.80105329516571e+006 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port6_port2_p2 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.13978752587401e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port6_port2_p3 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	5.33721279797821e+010 	3.88208408411310e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port6_port3_p1 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	2.16666961187778e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port6_port3_p2 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	1.38148736428337e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port6_port3_p3 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	-1.75646416707469e+010 	1.50395977768986e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port6_port4_p1 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.96964053709550e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port6_port4_p2 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.88462510318307e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port6_port4_p3 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	9.57369477165946e+010 	3.22486483351622e+010 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port6_port5_p1 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	3.74108139465422e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port6_port5_p2 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	2.92153191949078e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port6_port5_p3 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	-4.74723615989712e+010 	-8.54982158167148e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010
G_POLE_port6_port6_p1 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-4.14854779789202e+007 / 1.0 	3.92613467538825e+009 , 0.0
G_POLE_port6_port6_p2 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.75585631946697e+009 / 1.0 	5.13513753320332e+010 , 0.0
G_POLE_port6_port6_p3 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.65123498189666e+010 	-3.28428435379864e+011 , 0.0 / 1.0 	1.55180148415796e+011 , -2.41427481601416e+010


.ENDS  bbspice_subckt
***************************************


***************************************
* S-based subckt

 
*bbspice subcircuit with external port numbers.

*.SUBCKT bbspice_Case2_1mm		1 	2 	3 	4 	5 	6 	0 
*
*x_ 	1 	2 	3 	4 	5 	6 	0 	bbspice_Case2_1mm_subckt
*
*.ENDS  bbspice_Case2_1mm
***************************************
*.ENDL
