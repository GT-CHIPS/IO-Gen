
.PARAM tclk=1n l_tr=0.7m
