
.subckt IO_TX_ESD A VDDIO VSSIO
.ends
.subckt IO_RX_ESD A VDDIO VSSIO
.ends
