* Momentum eesofbbs_64 12.00 (*) built: Jan 14 2016
**************************************************
*.LIB Case4_1mm

*bbspice subcircuit with consecutive port numbers.

.SUBCKT bbspice_subckt	  port_1  port_2  port_3  port_4  port_5  port_6  gnd_0

* PORT_1
vi_1	port_1	_net_1	0.00000000000000e+000
vb_1	_net_4	_net_5	0.00000000000000e+000
R_Z0_1 	_net_1 	_net_2 	5.00000000000000e+001	NOISE=0
H_b_1	_net_2	gnd_0	vb_1	1.41421356237310e+001
E_v_1	_net_3	gnd_0	port_1	gnd_0	7.07106781186548e-002
H_i_1	_net_4	_net_3	vi_1	3.53553390593274e+000


G_POLE_port1_port1_p1 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-4.07455818618072e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port1_port1_p2 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.38246656805634e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port1_port1_p3 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.27672155296633e+010 	-2.46789224040305e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port1_port2_p1 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	3.67722415926790e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port1_port2_p2 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	2.32713817901723e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port1_port2_p3 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	-4.07624636294032e+010 	-1.14998115177392e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port1_port3_p1 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.08479094156762e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port1_port3_p2 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.41921658232922e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port1_port3_p3 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	1.03416516512980e+011 	2.86499874935292e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port1_port4_p1 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	2.23605629768335e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port1_port4_p2 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	1.01800131739065e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port1_port4_p3 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.48078044781903e+010 	1.72509936363303e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port1_port5_p1 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	4.24234821610131e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port1_port5_p2 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	-7.30263230766125e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port1_port5_p3 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	5.85492806425894e+010 	3.20229118148222e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port1_port6_p1 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	-4.79675394075645e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port1_port6_p2 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	7.84367252997538e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port1_port6_p3 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-2.94555712000663e+009 	6.55363538351850e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010

* PORT_2
vi_2	port_2	_net_6	0.00000000000000e+000
vb_2	_net_9	_net_10	0.00000000000000e+000
R_Z0_2 	_net_6 	_net_7 	5.00000000000000e+001	NOISE=0
H_b_2	_net_7	gnd_0	vb_2	1.41421356237310e+001
E_v_2	_net_8	gnd_0	port_2	gnd_0	7.07106781186548e-002
H_i_2	_net_9	_net_8	vi_2	3.53553390593274e+000


G_POLE_port2_port1_p1 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	3.67722415926790e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port2_port1_p2 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	2.32713817901723e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port2_port1_p3 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	-4.07624636294032e+010 	-1.14998115177392e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port2_port2_p1 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-4.12041613936215e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port2_port2_p2 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.32274713414487e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port2_port2_p3 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.21762543502408e+010 	-2.50643441247144e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port2_port3_p1 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	2.24117941016697e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port2_port3_p2 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	1.00975183655073e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port2_port3_p3 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	-1.49176054975383e+010 	1.70674384942834e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port2_port4_p1 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.03399134195575e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port2_port4_p2 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.47961016070037e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port2_port4_p3 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	1.02714777329723e+011 	2.94439174052776e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port2_port5_p1 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	-4.75939146846667e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port2_port5_p2 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	7.78068224244550e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port2_port5_p3 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-3.02949602376099e+009 	6.35098216547604e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port2_port6_p1 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	4.78688592297327e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port2_port6_p2 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	-7.91198270031207e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port2_port6_p3 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	5.78547655171478e+010 	3.34905642305741e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010

* PORT_3
vi_3	port_3	_net_11	0.00000000000000e+000
vb_3	_net_14	_net_15	0.00000000000000e+000
R_Z0_3 	_net_11 	_net_12 	5.00000000000000e+001	NOISE=0
H_b_3	_net_12	gnd_0	vb_3	1.41421356237310e+001
E_v_3	_net_13	gnd_0	port_3	gnd_0	7.07106781186548e-002
H_i_3	_net_14	_net_13	vi_3	3.53553390593274e+000


G_POLE_port3_port1_p1 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.08479094156762e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port3_port1_p2 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.41921658232922e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port3_port1_p3 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	1.03416516512980e+011 	2.86499874935292e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port3_port2_p1 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	2.24117941016697e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port3_port2_p2 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	1.00975183655073e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port3_port2_p3 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.49176054975383e+010 	1.70674384942834e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port3_port3_p1 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-5.08165468752521e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port3_port3_p2 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.04046719059154e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port3_port3_p3 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	-7.37118840126602e+008 	-8.62424978648745e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port3_port4_p1 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	4.60855567577912e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port3_port4_p2 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	3.14413374389205e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port3_port4_p3 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	-3.61290481099198e+010 	-1.27249921728204e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port3_port5_p1 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-2.06779085866474e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port3_port5_p2 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.40619433566568e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port3_port5_p3 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	1.03319728218245e+011 	2.85332782570241e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port3_port6_p1 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	2.20243188092829e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port3_port6_p2 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	1.04002112695715e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port3_port6_p3 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.53135413405720e+010 	1.68179354095860e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010

* PORT_4
vi_4	port_4	_net_16	0.00000000000000e+000
vb_4	_net_19	_net_20	0.00000000000000e+000
R_Z0_4 	_net_16 	_net_17 	5.00000000000000e+001	NOISE=0
H_b_4	_net_17	gnd_0	vb_4	1.41421356237310e+001
E_v_4	_net_18	gnd_0	port_4	gnd_0	7.07106781186548e-002
H_i_4	_net_19	_net_18	vi_4	3.53553390593274e+000


G_POLE_port4_port1_p1 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	2.23605629768335e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port4_port1_p2 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	1.01800131739065e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port4_port1_p3 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.48078044781903e+010 	1.72509936363303e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port4_port2_p1 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-2.03399134195575e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port4_port2_p2 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.47961016070037e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port4_port2_p3 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	1.02714777329723e+011 	2.94439174052776e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port4_port3_p1 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	4.60855567577912e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port4_port3_p2 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	3.14413374389205e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port4_port3_p3 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	-3.61290481099198e+010 	-1.27249921728204e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port4_port4_p1 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-5.03655559307382e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port4_port4_p2 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.09778294951803e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port4_port4_p3 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.41913788812858e+009 	-4.52084939539906e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port4_port5_p1 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	2.20575436038552e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port4_port5_p2 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	1.03521095093610e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port4_port5_p3 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.53572571023974e+010 	1.67376720126377e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port4_port6_p1 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-2.01668943905395e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port4_port6_p2 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.46869466910023e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port4_port6_p3 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	1.02604006569768e+011 	2.93516539705331e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010

* PORT_5
vi_5	port_5	_net_21	0.00000000000000e+000
vb_5	_net_24	_net_25	0.00000000000000e+000
R_Z0_5 	_net_21 	_net_22 	5.00000000000000e+001	NOISE=0
H_b_5	_net_22	gnd_0	vb_5	1.41421356237310e+001
E_v_5	_net_23	gnd_0	port_5	gnd_0	7.07106781186548e-002
H_i_5	_net_24	_net_23	vi_5	3.53553390593274e+000


G_POLE_port5_port1_p1 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	4.24234821610131e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port5_port1_p2 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	-7.30263230766125e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port5_port1_p3 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	5.85492806425894e+010 	3.20229118148222e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port5_port2_p1 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	-4.75939146846667e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port5_port2_p2 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	7.78068224244550e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port5_port2_p3 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-3.02949602376099e+009 	6.35098216547604e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port5_port3_p1 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.06779085866474e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port5_port3_p2 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.40619433566568e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port5_port3_p3 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	1.03319728218245e+011 	2.85332782570241e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port5_port4_p1 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	2.20575436038552e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port5_port4_p2 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	1.03521095093610e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port5_port4_p3 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.53572571023974e+010 	1.67376720126377e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port5_port5_p1 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-4.07005264028772e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port5_port5_p2 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.37539737880134e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port5_port5_p3 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.92280776029253e+010 	-2.91785805483410e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port5_port6_p1 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	3.67917597102580e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port5_port6_p2 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	2.30185267923358e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port5_port6_p3 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	-3.98558934894087e+010 	-1.17679413376158e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010

* PORT_6
vi_6	port_6	_net_26	0.00000000000000e+000
vb_6	_net_29	_net_30	0.00000000000000e+000
R_Z0_6 	_net_26 	_net_27 	5.00000000000000e+001	NOISE=0
H_b_6	_net_27	gnd_0	vb_6	1.41421356237310e+001
E_v_6	_net_28	gnd_0	port_6	gnd_0	7.07106781186548e-002
H_i_6	_net_29	_net_28	vi_6	3.53553390593274e+000


G_POLE_port6_port1_p1 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	-4.79675394075645e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port6_port1_p2 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	7.84367252997538e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port6_port1_p3 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.94555712000663e+009 	6.55363538351850e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port6_port2_p1 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	4.78688592297327e+006 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port6_port2_p2 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	-7.91198270031207e+008 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port6_port2_p3 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	5.78547655171478e+010 	3.34905642305741e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port6_port3_p1 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	2.20243188092829e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port6_port3_p2 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	1.04002112695715e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port6_port3_p3 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	-1.53135413405720e+010 	1.68179354095860e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port6_port4_p1 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.01668943905395e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port6_port4_p2 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.46869466910023e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port6_port4_p3 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	1.02604006569768e+011 	2.93516539705331e+010 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port6_port5_p1 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	3.67917597102580e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port6_port5_p2 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	2.30185267923358e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port6_port5_p3 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	-3.98558934894087e+010 	-1.17679413376158e+012 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010
G_POLE_port6_port6_p1 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-4.07782557300507e+007 / 1.0 	4.04385979201143e+009 , 0.0
G_POLE_port6_port6_p2 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.38680900083779e+009 / 1.0 	5.07786301984572e+010 , 0.0
G_POLE_port6_port6_p3 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.94621193941408e+010 	-2.88969958311878e+011 , 0.0 / 1.0 	1.65908975699895e+011 , -2.56524748697934e+010


.ENDS  bbspice_subckt
***************************************


***************************************
* S-based subckt

 
*bbspice subcircuit with external port numbers.

*.SUBCKT bbspice_Case4_1mm		1 	2 	3 	4 	5 	6 	0 
*
*x_ 	1 	2 	3 	4 	5 	6 	0 	bbspice_Case4_1mm_subckt

*.ENDS  bbspice_Case4_1mm
***************************************
*.ENDL
