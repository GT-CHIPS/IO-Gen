* Momentum eesofbbs_64 12.00 (*) built: Jan 14 2016
**************************************************
*.LIB Case2_5mm
*
**bbspice subcircuit with consecutive port numbers.
*
.SUBCKT bbspice_subckt	  port_1  port_2  port_3  port_4  port_5  port_6  gnd_0

* PORT_1
vi_1	port_1	_net_1	0.00000000000000e+000
vb_1	_net_4	_net_5	0.00000000000000e+000
R_Z0_1 	_net_1 	_net_2 	5.00000000000000e+001	NOISE=0
H_b_1	_net_2	gnd_0	vb_1	1.41421356237310e+001
E_v_1	_net_3	gnd_0	port_1	gnd_0	7.07106781186548e-002
H_i_1	_net_4	_net_3	vi_1	3.53553390593274e+000


G_POLE_port1_port1_p1 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-5.16376647440025e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port1_port1_p2 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-4.37677642412366e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port1_port1_p3 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	3.41802765937448e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port1_port1_p4 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	2.58533789020631e+007 	-1.68368266269750e+014 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port1_port1_p6 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	-3.73543824953017e+010 	-1.54650308595157e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port1_port2_p1 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	5.12909327868497e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port1_port2_p2 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	3.35258978028387e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port1_port2_p3 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	6.23805516296887e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port1_port2_p4 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.14614500952442e+011 	8.39420064284828e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port1_port2_p6 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	6.70067804803539e+010 	1.48137853497280e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port1_port3_p1 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.48775234790337e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port1_port3_p2 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.20692141237176e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port1_port3_p3 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-4.27910570349463e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port1_port3_p4 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	-7.71692856833600e+010 	7.41289287671111e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port1_port3_p6 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	1.82624108951087e+011 	2.08029317264670e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port1_port4_p1 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	2.50167084450331e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port1_port4_p2 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	2.22853716065277e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port1_port4_p3 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.50482942367729e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port1_port4_p4 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	-3.75530160023188e+010 	1.57365847239726e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port1_port4_p6 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	5.22875444002258e+010 	4.68277867220274e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port1_port5_p1 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	6.53170792868356e+006 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port1_port5_p2 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	1.77844103918858e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port1_port5_p3 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	-2.37126198765144e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port1_port5_p4 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	-5.70223568317921e+010 	2.82271143215208e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port1_port5_p6 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	1.39726879300353e+011 	1.23728298370728e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port1_port6_p1 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.21722994654052e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port1_port6_p2 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	1.29376854114771e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port1_port6_p3 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.34228553523945e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port1_port6_p4 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.69242620412669e+010 	-6.68766922377338e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port1_port6_p6 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	4.59705004479850e+010 	5.63210828908376e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010

* PORT_2
vi_2	port_2	_net_6	0.00000000000000e+000
vb_2	_net_9	_net_10	0.00000000000000e+000
R_Z0_2 	_net_6 	_net_7 	5.00000000000000e+001	NOISE=0
H_b_2	_net_7	gnd_0	vb_2	1.41421356237310e+001
E_v_2	_net_8	gnd_0	port_2	gnd_0	7.07106781186548e-002
H_i_2	_net_9	_net_8	vi_2	3.53553390593274e+000


G_POLE_port2_port1_p1 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	5.12909327868497e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port2_port1_p2 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	3.35258978028387e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port2_port1_p3 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	6.23805516296887e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port2_port1_p4 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.14614500952442e+011 	8.39420064284828e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port2_port1_p6 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	6.70067804803539e+010 	1.48137853497280e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port2_port2_p1 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-5.16944023186651e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port2_port2_p2 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-4.36057415562828e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port2_port2_p3 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	3.39751052293382e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port2_port2_p4 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.50949178681099e+009 	2.90934655565369e+012 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port2_port2_p6 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	-3.52257163642892e+010 	-2.19310821304026e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port2_port3_p1 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	2.49966634008121e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port2_port3_p2 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	2.23790374997684e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port2_port3_p3 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.50586765909324e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port2_port3_p4 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	-3.75815980069611e+010 	1.57002435502356e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port2_port3_p6 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	5.24038401338939e+010 	4.66901924157792e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port2_port4_p1 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.49413592674731e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port2_port4_p2 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.19060933370478e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port2_port4_p3 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-4.29378792277983e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port2_port4_p4 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	-7.80014395880595e+010 	7.38631632525658e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port2_port4_p6 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	1.83819186567992e+011 	2.07601156523263e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port2_port5_p1 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.22048412259134e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port2_port5_p2 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	1.30452152878455e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port2_port5_p3 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.34499417145498e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port2_port5_p4 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.70257985448857e+010 	-6.63685148607323e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port2_port5_p6 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	4.61825712289166e+010 	5.64254614490273e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port2_port6_p1 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	6.48879183406642e+006 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port2_port6_p2 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	1.78989419653635e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port2_port6_p3 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	-2.37812145411791e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port2_port6_p4 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	-5.76111737018675e+010 	2.82175481037578e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port2_port6_p6 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	1.40632412622813e+011 	1.23440735830423e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010

* PORT_3
vi_3	port_3	_net_11	0.00000000000000e+000
vb_3	_net_14	_net_15	0.00000000000000e+000
R_Z0_3 	_net_11 	_net_12 	5.00000000000000e+001	NOISE=0
H_b_3	_net_12	gnd_0	vb_3	1.41421356237310e+001
E_v_3	_net_13	gnd_0	port_3	gnd_0	7.07106781186548e-002
H_i_3	_net_14	_net_13	vi_3	3.53553390593274e+000


G_POLE_port3_port1_p1 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.48775234790337e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port3_port1_p2 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.20692141237176e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port3_port1_p3 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-4.27910570349463e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port3_port1_p4 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	-7.71692856833600e+010 	7.41289287671111e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port3_port1_p6 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	1.82624108951087e+011 	2.08029317264670e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port3_port2_p1 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	2.49966634008121e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port3_port2_p2 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	2.23790374997684e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port3_port2_p3 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	-2.50586765909324e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port3_port2_p4 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	-3.75815980069611e+010 	1.57002435502356e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port3_port2_p6 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	5.24038401338939e+010 	4.66901924157792e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port3_port3_p1 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-6.91420906804675e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port3_port3_p2 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-4.33732323758211e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port3_port3_p3 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	2.61307688195182e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port3_port3_p4 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	-2.49876423788303e+010 	1.88391650477857e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port3_port3_p6 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	1.98990216370140e+010 	2.86117763977907e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port3_port4_p1 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	6.33261844898431e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port3_port4_p2 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	6.08230684652888e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port3_port4_p3 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	6.42161476615777e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port3_port4_p4 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.18627107591160e+011 	6.27071114972499e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port3_port4_p6 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	9.21543992845832e+010 	3.56974657642511e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port3_port5_p1 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-2.48235870250039e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port3_port5_p2 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-2.24741586332042e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port3_port5_p3 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-4.28095704168651e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port3_port5_p4 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	-7.74334837830134e+010 	7.34986833501100e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port3_port5_p6 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	1.83435513823176e+011 	2.06826568352413e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port3_port6_p1 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	2.51008538245484e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port3_port6_p2 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	2.19759197476460e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port3_port6_p3 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	-2.51399709891963e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port3_port6_p4 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	-3.79590298997676e+010 	1.55509334983728e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port3_port6_p6 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	5.30734135327590e+010 	4.62039608707928e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010

* PORT_4
vi_4	port_4	_net_16	0.00000000000000e+000
vb_4	_net_19	_net_20	0.00000000000000e+000
R_Z0_4 	_net_16 	_net_17 	5.00000000000000e+001	NOISE=0
H_b_4	_net_17	gnd_0	vb_4	1.41421356237310e+001
E_v_4	_net_18	gnd_0	port_4	gnd_0	7.07106781186548e-002
H_i_4	_net_19	_net_18	vi_4	3.53553390593274e+000


G_POLE_port4_port1_p1 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	2.50167084450331e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port4_port1_p2 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	2.22853716065277e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port4_port1_p3 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.50482942367729e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port4_port1_p4 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	-3.75530160023188e+010 	1.57365847239726e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port4_port1_p6 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	5.22875444002258e+010 	4.68277867220274e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port4_port2_p1 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-2.49413592674731e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port4_port2_p2 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-2.19060933370478e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port4_port2_p3 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-4.29378792277983e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port4_port2_p4 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	-7.80014395880595e+010 	7.38631632525658e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port4_port2_p6 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	1.83819186567992e+011 	2.07601156523263e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port4_port3_p1 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	6.33261844898431e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port4_port3_p2 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	6.08230684652888e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port4_port3_p3 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	6.42161476615777e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port4_port3_p4 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	-1.18627107591160e+011 	6.27071114972499e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port4_port3_p6 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	9.21543992845832e+010 	3.56974657642511e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port4_port4_p1 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-6.92194512476123e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port4_port4_p2 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-4.31150403938375e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port4_port4_p3 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	2.58904573567651e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port4_port4_p4 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	-2.62320489617449e+010 	1.82080540919723e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port4_port4_p6 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	2.16233618546115e+010 	2.76355057701512e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port4_port5_p1 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	2.50732315611353e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port4_port5_p2 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	2.20639333849459e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port4_port5_p3 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	-2.51714237226766e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port4_port5_p4 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	-3.80101795118432e+010 	1.55638325913989e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port4_port5_p6 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	5.31238021154403e+010 	4.62450871760780e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port4_port6_p1 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-2.49025474947673e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port4_port6_p2 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-2.22030919242913e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port4_port6_p3 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-4.29980835855646e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port4_port6_p4 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	-7.83653898925980e+010 	7.33677160030575e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port4_port6_p6 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	1.84782964126266e+011 	2.06564164910946e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010

* PORT_5
vi_5	port_5	_net_21	0.00000000000000e+000
vb_5	_net_24	_net_25	0.00000000000000e+000
R_Z0_5 	_net_21 	_net_22 	5.00000000000000e+001	NOISE=0
H_b_5	_net_22	gnd_0	vb_5	1.41421356237310e+001
E_v_5	_net_23	gnd_0	port_5	gnd_0	7.07106781186548e-002
H_i_5	_net_24	_net_23	vi_5	3.53553390593274e+000


G_POLE_port5_port1_p1 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	6.53170792868356e+006 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port5_port1_p2 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	1.77844103918858e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port5_port1_p3 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.37126198765144e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port5_port1_p4 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	-5.70223568317921e+010 	2.82271143215208e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port5_port1_p6 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	1.39726879300353e+011 	1.23728298370728e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port5_port2_p1 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.22048412259134e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port5_port2_p2 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	1.30452152878455e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port5_port2_p3 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.34499417145498e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port5_port2_p4 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.70257985448857e+010 	-6.63685148607323e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port5_port2_p6 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	4.61825712289166e+010 	5.64254614490273e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port5_port3_p1 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.48235870250039e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port5_port3_p2 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.24741586332042e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port5_port3_p3 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-4.28095704168651e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port5_port3_p4 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	-7.74334837830134e+010 	7.34986833501100e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port5_port3_p6 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	1.83435513823176e+011 	2.06826568352413e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port5_port4_p1 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	2.50732315611353e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port5_port4_p2 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	2.20639333849459e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port5_port4_p3 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.51714237226766e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port5_port4_p4 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	-3.80101795118432e+010 	1.55638325913989e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port5_port4_p6 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	5.31238021154403e+010 	4.62450871760780e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port5_port5_p1 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-5.17389708871582e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port5_port5_p2 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-4.35959338528708e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port5_port5_p3 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	3.45118944813846e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port5_port5_p4 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	-3.05844802826569e+008 	1.39795545970692e+013 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port5_port5_p6 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	-3.62946816363379e+010 	-6.11212792277594e+009 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port5_port6_p1 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	5.13503939459400e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port5_port6_p2 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	3.34462778421159e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port5_port6_p3 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	6.26947434600147e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port5_port6_p4 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.14527902031426e+011 	8.29381696050805e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port5_port6_p6 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	6.76926167568361e+010 	1.40010683334729e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010

* PORT_6
vi_6	port_6	_net_26	0.00000000000000e+000
vb_6	_net_29	_net_30	0.00000000000000e+000
R_Z0_6 	_net_26 	_net_27 	5.00000000000000e+001	NOISE=0
H_b_6	_net_27	gnd_0	vb_6	1.41421356237310e+001
E_v_6	_net_28	gnd_0	port_6	gnd_0	7.07106781186548e-002
H_i_6	_net_29	_net_28	vi_6	3.53553390593274e+000


G_POLE_port6_port1_p1 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.21722994654052e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port6_port1_p2 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	1.29376854114771e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port6_port1_p3 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.34228553523945e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port6_port1_p4 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.69242620412669e+010 	-6.68766922377338e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port6_port1_p6 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	4.59705004479850e+010 	5.63210828908376e+010 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port6_port2_p1 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	6.48879183406642e+006 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port6_port2_p2 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	1.78989419653635e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port6_port2_p3 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	-2.37812145411791e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port6_port2_p4 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	-5.76111737018675e+010 	2.82175481037578e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port6_port2_p6 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	1.40632412622813e+011 	1.23440735830423e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port6_port3_p1 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	2.51008538245484e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port6_port3_p2 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	2.19759197476460e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port6_port3_p3 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.51399709891963e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port6_port3_p4 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	-3.79590298997676e+010 	1.55509334983728e+011 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port6_port3_p6 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	5.30734135327590e+010 	4.62039608707928e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port6_port4_p1 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.49025474947673e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port6_port4_p2 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.22030919242913e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port6_port4_p3 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-4.29980835855646e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port6_port4_p4 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	-7.83653898925980e+010 	7.33677160030575e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port6_port4_p6 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	1.84782964126266e+011 	2.06564164910946e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port6_port5_p1 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	5.13503939459400e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port6_port5_p2 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	3.34462778421159e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port6_port5_p3 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	6.26947434600147e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port6_port5_p4 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.14527902031426e+011 	8.29381696050805e+010 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port6_port5_p6 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	6.76926167568361e+010 	1.40010683334729e+011 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010
G_POLE_port6_port6_p1 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-5.17972340200316e+007 / 1.0 	2.34061526025922e+009 , 0.0
G_POLE_port6_port6_p2 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-4.34503522818358e+008 / 1.0 	1.48610484404771e+010 , 0.0
G_POLE_port6_port6_p3 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	3.44230804950835e+010 / 1.0 	5.33129796941333e+010 , 0.0
G_POLE_port6_port6_p4 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.75280157070113e+009 	2.45320431843880e+012 , 0.0 / 1.0 	5.76988198652384e+010 , -1.46428062934995e+010
G_POLE_port6_port6_p6 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	-3.35589158609996e+010 	-9.62370452472592e+009 , 0.0 / 1.0 	1.44608877342323e+011 , -1.30788559350683e+010


.ENDS  bbspice_subckt
***************************************


***************************************
* S-based subckt

 
*bbspice subcircuit with external port numbers.

*.SUBCKT bbspice_Case2_5mm		1 	2 	3 	4 	5 	6 	0 
*
*x_ 	1 	2 	3 	4 	5 	6 	0 	bbspice_Case2_5mm_subckt
*
*.ENDS  bbspice_Case2_5mm
****************************************
*.ENDL
