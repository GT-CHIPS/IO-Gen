* Momentum eesofbbs_64 12.00 (*) built: Jan 14 2016
**************************************************
*.LIB Case1_1mm

*bbspice subcircuit with consecutive port numbers.

.SUBCKT bbspice_subckt	  port_1  port_2  port_3  port_4  port_5  port_6  gnd_0

* PORT_1
vi_1	port_1	_net_1	0.00000000000000e+000
vb_1	_net_4	_net_5	0.00000000000000e+000
R_Z0_1 	_net_1 	_net_2 	5.00000000000000e+001	NOISE=0
H_b_1	_net_2	gnd_0	vb_1	1.41421356237310e+001
E_v_1	_net_3	gnd_0	port_1	gnd_0	7.07106781186548e-002
H_i_1	_net_4	_net_3	vi_1	3.53553390593274e+000


G_POLE_port1_port1_p1 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-5.33560622331382e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port1_port1_p2 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-8.31355881272227e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port1_port1_p3 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	6.30666155524492e+010 	2.16447063846186e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port1_port2_p1 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	5.29544409527549e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port1_port2_p2 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	-3.48590627139831e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port1_port2_p3 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	1.07919683267886e+011 	2.36713712186771e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port1_port3_p1 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.26692547784000e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port1_port3_p2 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	3.06711520655744e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port1_port3_p3 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	1.40158095860273e+010 	-2.72038849901249e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port1_port4_p1 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	1.49679133484342e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port1_port4_p2 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	-6.26377555159599e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port1_port4_p3 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	5.35816483843443e+009 	-4.81072184602690e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port1_port5_p1 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	3.58736982235008e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port1_port5_p2 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	1.80119366487210e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port1_port5_p3 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	-2.26872342410485e+010 	7.52095700049337e+010 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port1_port6_p1 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	-3.00804559016111e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port1_port6_p2 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	4.31393678051842e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port1_port6_p3 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.47909241908385e+010 	2.08198425060769e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010

* PORT_2
vi_2	port_2	_net_6	0.00000000000000e+000
vb_2	_net_9	_net_10	0.00000000000000e+000
R_Z0_2 	_net_6 	_net_7 	5.00000000000000e+001	NOISE=0
H_b_2	_net_7	gnd_0	vb_2	1.41421356237310e+001
E_v_2	_net_8	gnd_0	port_2	gnd_0	7.07106781186548e-002
H_i_2	_net_9	_net_8	vi_2	3.53553390593274e+000


G_POLE_port2_port1_p1 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	5.29544409527549e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port2_port1_p2 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	-3.48590627139831e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port2_port1_p3 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	1.07919683267886e+011 	2.36713712186771e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port2_port2_p1 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-5.37907075518587e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port2_port2_p2 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.93579148483421e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port2_port2_p3 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	6.46563106635028e+010 	2.14804089379388e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port2_port3_p1 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	1.49840846342941e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port2_port3_p2 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	-6.23155706257594e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port2_port3_p3 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	5.39774650508564e+009 	-4.77694363576609e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port2_port4_p1 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.26636486923826e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port2_port4_p2 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	3.07887566657017e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port2_port4_p3 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	1.40295984953044e+010 	-2.73549155830517e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port2_port5_p1 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	-3.00161981054639e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port2_port5_p2 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	4.34726768343767e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port2_port5_p3 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.48108229619285e+010 	2.08433475342320e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port2_port6_p1 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	3.60689654635913e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port2_port6_p2 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	1.82720211908661e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port2_port6_p3 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	-2.32345689906528e+010 	7.58892810998858e+010 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010

* PORT_3
vi_3	port_3	_net_11	0.00000000000000e+000
vb_3	_net_14	_net_15	0.00000000000000e+000
R_Z0_3 	_net_11 	_net_12 	5.00000000000000e+001	NOISE=0
H_b_3	_net_12	gnd_0	vb_3	1.41421356237310e+001
E_v_3	_net_13	gnd_0	port_3	gnd_0	7.07106781186548e-002
H_i_3	_net_14	_net_13	vi_3	3.53553390593274e+000


G_POLE_port3_port1_p1 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.26692547784000e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port3_port1_p2 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	3.06711520655744e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port3_port1_p3 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	1.40158095860273e+010 	-2.72038849901249e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port3_port2_p1 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	1.49840846342941e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port3_port2_p2 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	-6.23155706257594e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port3_port2_p3 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	5.39774650508564e+009 	-4.77694363576609e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port3_port3_p1 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.82662725091519e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port3_port3_p2 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	7.38142602498057e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port3_port3_p3 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	5.96851766419431e+010 	1.88078544184086e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port3_port4_p1 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	4.90569265319912e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port3_port4_p2 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	-2.81853078257026e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port3_port4_p3 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	1.02569816709294e+011 	2.40893776280294e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port3_port5_p1 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.21561741720461e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port3_port5_p2 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	3.04605418703101e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port3_port5_p3 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	1.39122188958931e+010 	-2.71203749150642e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port3_port6_p1 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	1.44451682762622e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port3_port6_p2 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	-5.17925823012218e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port3_port6_p3 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	4.61886479031634e+009 	-5.61971867606867e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010

* PORT_4
vi_4	port_4	_net_16	0.00000000000000e+000
vb_4	_net_19	_net_20	0.00000000000000e+000
R_Z0_4 	_net_16 	_net_17 	5.00000000000000e+001	NOISE=0
H_b_4	_net_17	gnd_0	vb_4	1.41421356237310e+001
E_v_4	_net_18	gnd_0	port_4	gnd_0	7.07106781186548e-002
H_i_4	_net_19	_net_18	vi_4	3.53553390593274e+000


G_POLE_port4_port1_p1 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	1.49679133484342e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port4_port1_p2 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	-6.26377555159599e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port4_port1_p3 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	5.35816483843443e+009 	-4.81072184602690e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port4_port2_p1 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.26636486923826e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port4_port2_p2 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	3.07887566657017e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port4_port2_p3 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	1.40295984953044e+010 	-2.73549155830517e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port4_port3_p1 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	4.90569265319912e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port4_port3_p2 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	-2.81853078257026e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port4_port3_p3 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	1.02569816709294e+011 	2.40893776280294e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port4_port4_p1 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.84031123186208e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port4_port4_p2 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	6.61603709195879e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port4_port4_p3 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	6.07680258216784e+010 	1.87416497768289e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port4_port5_p1 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	1.45869821788867e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port4_port5_p2 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	-4.32601177769690e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port4_port5_p3 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	4.45788568106607e+009 	-5.86614120895877e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port4_port6_p1 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.22765422177869e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port4_port6_p2 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	3.09718962541711e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port4_port6_p3 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	1.32151603198636e+010 	-2.93623313308497e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010

* PORT_5
vi_5	port_5	_net_21	0.00000000000000e+000
vb_5	_net_24	_net_25	0.00000000000000e+000
R_Z0_5 	_net_21 	_net_22 	5.00000000000000e+001	NOISE=0
H_b_5	_net_22	gnd_0	vb_5	1.41421356237310e+001
E_v_5	_net_23	gnd_0	port_5	gnd_0	7.07106781186548e-002
H_i_5	_net_24	_net_23	vi_5	3.53553390593274e+000


G_POLE_port5_port1_p1 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	3.58736982235008e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port5_port1_p2 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	1.80119366487210e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port5_port1_p3 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.26872342410485e+010 	7.52095700049337e+010 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port5_port2_p1 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	-3.00161981054639e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port5_port2_p2 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	4.34726768343767e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port5_port2_p3 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.48108229619285e+010 	2.08433475342320e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port5_port3_p1 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.21561741720461e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port5_port3_p2 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	3.04605418703101e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port5_port3_p3 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	1.39122188958931e+010 	-2.71203749150642e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port5_port4_p1 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	1.45869821788867e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port5_port4_p2 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	-4.32601177769690e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port5_port4_p3 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	4.45788568106607e+009 	-5.86614120895877e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port5_port5_p1 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-5.31315973330213e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port5_port5_p2 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.53017879576446e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port5_port5_p3 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	6.54961405493644e+010 	2.10649148356943e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port5_port6_p1 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	5.29430135367236e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port5_port6_p2 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	-3.51013300885023e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port5_port6_p3 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	1.09154338789540e+011 	2.34504145289623e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010

* PORT_6
vi_6	port_6	_net_26	0.00000000000000e+000
vb_6	_net_29	_net_30	0.00000000000000e+000
R_Z0_6 	_net_26 	_net_27 	5.00000000000000e+001	NOISE=0
H_b_6	_net_27	gnd_0	vb_6	1.41421356237310e+001
E_v_6	_net_28	gnd_0	port_6	gnd_0	7.07106781186548e-002
H_i_6	_net_29	_net_28	vi_6	3.53553390593274e+000


G_POLE_port6_port1_p1 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	-3.00804559016111e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port6_port1_p2 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	4.31393678051842e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port6_port1_p3 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.47909241908385e+010 	2.08198425060769e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port6_port2_p1 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	3.60689654635913e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port6_port2_p2 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	1.82720211908661e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port6_port2_p3 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.32345689906528e+010 	7.58892810998858e+010 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port6_port3_p1 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	1.44451682762622e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port6_port3_p2 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	-5.17925823012218e+010 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port6_port3_p3 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	4.61886479031634e+009 	-5.61971867606867e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port6_port4_p1 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.22765422177869e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port6_port4_p2 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	3.09718962541711e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port6_port4_p3 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	1.32151603198636e+010 	-2.93623313308497e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port6_port5_p1 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	5.29430135367236e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port6_port5_p2 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	-3.51013300885023e+012 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port6_port5_p3 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	1.09154338789540e+011 	2.34504145289623e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010
G_POLE_port6_port6_p1 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-5.34783319324923e+008 / 1.0 	3.21249370645228e+010 , 0.0
G_POLE_port6_port6_p2 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.70403113448116e+011 / 1.0 	1.49374267959163e+013 , 0.0
G_POLE_port6_port6_p3 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	6.54506524428813e+010 	2.11406435223477e+011 , 0.0 / 1.0 	1.62736285787277e+011 , -1.14414366404791e+010


.ENDS  bbspice_subckt
***************************************


***************************************
* S-based subckt

 
*bbspice subcircuit with external port numbers.

*.SUBCKT bbspice_Case1_1mm		1 	2 	3 	4 	5 	6 	0 
*
*x_ 	1 	2 	3 	4 	5 	6 	0 	bbspice_Case1_1mm_subckt
*
*.ENDS  bbspice_Case1_1mm
****************************************
*.ENDL
