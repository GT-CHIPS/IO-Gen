* Momentum eesofbbs_64 12.00 (*) built: Jan 14 2016
**************************************************
*.LIB GSG_Case2_C4_5mmTLIN_C4_20GHz

*bbspice subcircuit with consecutive port numbers.

.SUBCKT bbspice_GSG_Case2_5mm_20GHz_subckt	  port_1  port_2  gnd_0

* PORT_1
vi_1	port_1	_net_1	0.00000000000000e+000
vb_1	_net_4	_net_5	0.00000000000000e+000
R_Z0_1 	_net_1 	_net_2 	5.00000000000000e+001	NOISE=0
H_b_1	_net_2	gnd_0	vb_1	1.41421356237310e+001
E_v_1	_net_3	gnd_0	port_1	gnd_0	7.07106781186548e-002
H_i_1	_net_4	_net_3	vi_1	3.53553390593274e+000


G_port1_port1 	_net_5	gnd_0	_net_5	gnd_0	3.29246449279721e-001
G_POLE_port1_port1_p1 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-8.95435158162820e+005 / 1.0 	8.43404417143702e+008 , 0.0
G_POLE_port1_port1_p2 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-4.13230067694628e+007 / 1.0 	2.38304952910240e+009 , 0.0
G_POLE_port1_port1_p3 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	7.24096498011585e+007 / 1.0 	4.50193013601027e+009 , 0.0
G_POLE_port1_port1_p4 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-5.16485403884426e+008 / 1.0 	9.56139413182203e+009 , 0.0
G_POLE_port1_port1_p5 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	1.08424464755049e+012 / 1.0 	9.95288743873958e+010 , 0.0
G_POLE_port1_port1_p6 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.28578568417364e+012 / 1.0 	1.16764351558112e+011 , 0.0
G_POLE_port1_port1_p7 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.00810941514175e+007 	-5.98147081729803e+009 , 0.0 / 1.0 	1.70137986630926e+009 , -8.40128737089965e+008
G_POLE_port1_port1_p9 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	3.84698891481663e+007 	-2.02472632530970e+009 , 0.0 / 1.0 	2.02411733488166e+009 , -8.79499553772000e+008
G_POLE_port1_port1_p11 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	3.28203811243767e+010 	-5.62601796852377e+009 , 0.0 / 1.0 	5.05577642516889e+010 , -5.36604122710960e+009
G_POLE_port1_port1_p13 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	2.17133976279853e+009 	5.79460214762948e+011 , 0.0 / 1.0 	3.91666816946069e+010 , -1.33316672667639e+010
G_POLE_port1_port1_p15 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	-4.18248338979271e+009 	-2.76214029249272e+010 , 0.0 / 1.0 	4.31674556130857e+010 , -1.71645028512267e+010
G_POLE_port1_port1_p17 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	9.11886060717353e+010 	8.39731439077971e+009 , 0.0 / 1.0 	6.42548226679118e+010 , -1.99085423767346e+010
G_POLE_port1_port2_p1 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	3.16417941291129e+006 / 1.0 	8.43404417143702e+008 , 0.0
G_POLE_port1_port2_p2 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.88256366729719e+007 / 1.0 	2.38304952910240e+009 , 0.0
G_POLE_port1_port2_p3 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	2.65285645121548e+008 / 1.0 	4.50193013601027e+009 , 0.0
G_POLE_port1_port2_p4 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	-2.81313331024437e+008 / 1.0 	9.56139413182203e+009 , 0.0
G_POLE_port1_port2_p5 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	1.39404336181841e+012 / 1.0 	9.95288743873958e+010 , 0.0
G_POLE_port1_port2_p6 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.34944437135900e+012 / 1.0 	1.16764351558112e+011 , 0.0
G_POLE_port1_port2_p7 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.05618449322348e+006 	-1.90815937472521e+011 , 0.0 / 1.0 	1.70137986630926e+009 , -8.40128737089965e+008
G_POLE_port1_port2_p9 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	3.78735654988831e+007 	-1.32894778468689e+010 , 0.0 / 1.0 	2.02411733488166e+009 , -8.79499553772000e+008
G_POLE_port1_port2_p11 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	2.25242772146298e+009 	-7.37016887507343e+011 , 0.0 / 1.0 	5.05577642516889e+010 , -5.36604122710960e+009
G_POLE_port1_port2_p13 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.27562005358579e+009 	-6.67118889421912e+011 , 0.0 / 1.0 	3.91666816946069e+010 , -1.33316672667639e+010
G_POLE_port1_port2_p15 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	5.19457447553975e+010 	8.71323623248519e+010 , 0.0 / 1.0 	4.31674556130857e+010 , -1.71645028512267e+010
G_POLE_port1_port2_p17 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	-7.42352485284662e+010 	4.68903885673835e+011 , 0.0 / 1.0 	6.42548226679118e+010 , -1.99085423767346e+010

* PORT_2
vi_2	port_2	_net_6	0.00000000000000e+000
vb_2	_net_9	_net_10	0.00000000000000e+000
R_Z0_2 	_net_6 	_net_7 	5.00000000000000e+001	NOISE=0
H_b_2	_net_7	gnd_0	vb_2	1.41421356237310e+001
E_v_2	_net_8	gnd_0	port_2	gnd_0	7.07106781186548e-002
H_i_2	_net_9	_net_8	vi_2	3.53553390593274e+000


G_POLE_port2_port1_p1 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	3.16417941291129e+006 / 1.0 	8.43404417143702e+008 , 0.0
G_POLE_port2_port1_p2 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.88256366729719e+007 / 1.0 	2.38304952910240e+009 , 0.0
G_POLE_port2_port1_p3 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	2.65285645121548e+008 / 1.0 	4.50193013601027e+009 , 0.0
G_POLE_port2_port1_p4 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.81313331024437e+008 / 1.0 	9.56139413182203e+009 , 0.0
G_POLE_port2_port1_p5 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	1.39404336181841e+012 / 1.0 	9.95288743873958e+010 , 0.0
G_POLE_port2_port1_p6 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.34944437135900e+012 / 1.0 	1.16764351558112e+011 , 0.0
G_POLE_port2_port1_p7 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.05618449322348e+006 	-1.90815937472521e+011 , 0.0 / 1.0 	1.70137986630926e+009 , -8.40128737089965e+008
G_POLE_port2_port1_p9 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	3.78735654988831e+007 	-1.32894778468689e+010 , 0.0 / 1.0 	2.02411733488166e+009 , -8.79499553772000e+008
G_POLE_port2_port1_p11 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	2.25242772146298e+009 	-7.37016887507343e+011 , 0.0 / 1.0 	5.05577642516889e+010 , -5.36604122710960e+009
G_POLE_port2_port1_p13 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.27562005358579e+009 	-6.67118889421912e+011 , 0.0 / 1.0 	3.91666816946069e+010 , -1.33316672667639e+010
G_POLE_port2_port1_p15 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	5.19457447553975e+010 	8.71323623248519e+010 , 0.0 / 1.0 	4.31674556130857e+010 , -1.71645028512267e+010
G_POLE_port2_port1_p17 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	-7.42352485284662e+010 	4.68903885673835e+011 , 0.0 / 1.0 	6.42548226679118e+010 , -1.99085423767346e+010
G_port2_port2 	_net_10	gnd_0	_net_10	gnd_0	3.30682548466158e-001
G_POLE_port2_port2_p1 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-9.20782875111350e+005 / 1.0 	8.43404417143702e+008 , 0.0
G_POLE_port2_port2_p2 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-4.07718984060499e+007 / 1.0 	2.38304952910240e+009 , 0.0
G_POLE_port2_port2_p3 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	6.97590088471373e+007 / 1.0 	4.50193013601027e+009 , 0.0
G_POLE_port2_port2_p4 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-5.11587946530061e+008 / 1.0 	9.56139413182203e+009 , 0.0
G_POLE_port2_port2_p5 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	1.09443742859870e+012 / 1.0 	9.95288743873958e+010 , 0.0
G_POLE_port2_port2_p6 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.29800542330814e+012 / 1.0 	1.16764351558112e+011 , 0.0
G_POLE_port2_port2_p7 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.01886557399408e+007 	-5.80405260722360e+009 , 0.0 / 1.0 	1.70137986630926e+009 , -8.40128737089965e+008
G_POLE_port2_port2_p9 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	3.83031280149251e+007 	-1.93487548078757e+009 , 0.0 / 1.0 	2.02411733488166e+009 , -8.79499553772000e+008
G_POLE_port2_port2_p11 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	3.32851124401047e+010 	-5.13094164598547e+009 , 0.0 / 1.0 	5.05577642516889e+010 , -5.36604122710960e+009
G_POLE_port2_port2_p13 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	2.41177195778636e+009 	5.52043261326268e+011 , 0.0 / 1.0 	3.91666816946069e+010 , -1.33316672667639e+010
G_POLE_port2_port2_p15 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.67364635712772e+009 	-7.82976362005828e+010 , 0.0 / 1.0 	4.31674556130857e+010 , -1.71645028512267e+010
G_POLE_port2_port2_p17 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	9.06725922159162e+010 	4.39083098557743e+009 , 0.0 / 1.0 	6.42548226679118e+010 , -1.99085423767346e+010


.ENDS  bbspice_GSG_Case2_5mm_20GHz_subckt
***************************************


***************************************
* S-based subckt

 
*bbspice subcircuit with external port numbers.

*.SUBCKT bbspice_GSG_Case2_C4_5mmTLIN_C4_20GHz		1 	2 	0 
*
*x_ 	1 	2 	0 	bbspice_GSG_Case2_C4_5mmTLIN_C4_20GHz_subckt
*
*.ENDS  bbspice_GSG_Case2_C4_5mmTLIN_C4_20GHz
****************************************
*.ENDL
