* Momentum eesofbbs_64 12.00 (*) built: Jan 14 2016
**************************************************
*.LIB Case4_10mm

*bbspice subcircuit with consecutive port numbers.

.SUBCKT bbspice_subckt	  port_1  port_2  port_3  port_4  port_5  port_6  gnd_0

* PORT_1
vi_1	port_1	_net_1	0.00000000000000e+000
vb_1	_net_4	_net_5	0.00000000000000e+000
R_Z0_1 	_net_1 	_net_2 	5.00000000000000e+001	NOISE=0
H_b_1	_net_2	gnd_0	vb_1	1.41421356237310e+001
E_v_1	_net_3	gnd_0	port_1	gnd_0	7.07106781186548e-002
H_i_1	_net_4	_net_3	vi_1	3.53553390593274e+000


G_POLE_port1_port1_p1 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	-8.49294465899445e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port1_port1_p2 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0  	6.60392125524830e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port1_port1_p3 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	8.25151696822376e+009 	4.23141117802762e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port1_port1_p5 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.23145151664942e+010 	3.16113855305808e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port1_port1_p7 	_net_5 	gnd_0 	POLE 	_net_5 	gnd_0 	7.98655907321926e+008 	8.59191672164281e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port1_port2_p1 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	8.17552955909611e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port1_port2_p2 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.23500346794900e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port1_port2_p3 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	2.31520733441888e+010 	3.27311362389721e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port1_port2_p5 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	-6.25315049407953e+009 	-2.68223856277640e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port1_port2_p7 	_net_5 	gnd_0 	POLE 	_net_10 	gnd_0 	4.62969191443515e+009 	-5.98452665502175e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port1_port3_p1 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.65334497161625e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port1_port3_p2 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0  	3.72090655250536e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port1_port3_p3 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	-8.15745392526853e+008 	1.96340124318664e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port1_port3_p5 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	-4.01595725118987e+009 	-5.04466643655448e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port1_port3_p7 	_net_5 	gnd_0 	POLE 	_net_15 	gnd_0 	3.62923575837272e+009 	2.16260786971802e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port1_port4_p1 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	3.32048496878048e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port1_port4_p2 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.35988352969782e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port1_port4_p3 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	-3.29885451651886e+008 	3.69688277466882e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port1_port4_p5 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	-8.09091751240442e+009 	1.27427420869376e+009 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port1_port4_p7 	_net_5 	gnd_0 	POLE 	_net_20 	gnd_0 	8.14616163766072e+009 	6.65606949405473e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port1_port5_p1 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	2.38180432316301e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port1_port5_p2 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0  	2.39295455907431e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port1_port5_p3 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.05209892494071e+010 	2.57606540413510e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port1_port5_p5 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	-2.12431904104578e+009 	-2.11874964036513e+011 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port1_port5_p7 	_net_5 	gnd_0 	POLE 	_net_25 	gnd_0 	7.55015440369252e+009 	5.56028200209978e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port1_port6_p1 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	-2.14994539100996e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port1_port6_p2 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0  	1.34173277083232e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port1_port6_p3 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-9.22512997184087e+009 	2.82385839737405e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port1_port6_p5 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-2.78597977624556e+009 	-7.99222224234456e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port1_port6_p7 	_net_5 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.21459579971251e+009 	-5.14290952085335e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010

* PORT_2
vi_2	port_2	_net_6	0.00000000000000e+000
vb_2	_net_9	_net_10	0.00000000000000e+000
R_Z0_2 	_net_6 	_net_7 	5.00000000000000e+001	NOISE=0
H_b_2	_net_7	gnd_0	vb_2	1.41421356237310e+001
E_v_2	_net_8	gnd_0	port_2	gnd_0	7.07106781186548e-002
H_i_2	_net_9	_net_8	vi_2	3.53553390593274e+000


G_POLE_port2_port1_p1 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	8.17552955909611e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port2_port1_p2 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.23500346794900e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port2_port1_p3 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	2.31520733441888e+010 	3.27311362389721e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port2_port1_p5 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	-6.25315049407953e+009 	-2.68223856277640e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port2_port1_p7 	_net_10 	gnd_0 	POLE 	_net_5 	gnd_0 	4.62969191443515e+009 	-5.98452665502175e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port2_port2_p1 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	-8.54370235292667e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port2_port2_p2 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0  	6.29175997575996e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port2_port2_p3 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	8.19727112437419e+009 	4.24214740605918e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port2_port2_p5 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.23656048407824e+010 	3.01896496523912e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port2_port2_p7 	_net_10 	gnd_0 	POLE 	_net_10 	gnd_0 	6.12971230129083e+008 	1.07071491440602e+012 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port2_port3_p1 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	3.30221042406057e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port2_port3_p2 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.51357824300096e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port2_port3_p3 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	-3.83896395732270e+008 	3.19628057927558e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port2_port3_p5 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	-7.96718679484474e+009 	5.50498003374687e+008 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port2_port3_p7 	_net_10 	gnd_0 	POLE 	_net_15 	gnd_0 	8.21479656290914e+009 	6.50142918198976e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port2_port4_p1 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.65578509876181e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port2_port4_p2 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0  	3.76406180657276e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port2_port4_p3 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.08800100515845e+009 	1.52634465650035e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port2_port4_p5 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	-4.25729105076331e+009 	-4.79159323433055e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port2_port4_p7 	_net_10 	gnd_0 	POLE 	_net_20 	gnd_0 	3.71033331149815e+009 	2.94237264253304e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port2_port5_p1 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	-2.17049499682876e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port2_port5_p2 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0  	1.32455533654710e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port2_port5_p3 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-9.24479371195703e+009 	2.81748019695366e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port2_port5_p5 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-2.64409687181222e+009 	-8.61126622278852e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port2_port5_p7 	_net_10 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.16774917735257e+009 	-5.25465779412074e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port2_port6_p1 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	2.37875391275076e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port2_port6_p2 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0  	2.43560461434402e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port2_port6_p3 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.08290404440687e+010 	2.55973078442315e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port2_port6_p5 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	-2.23526944528328e+009 	-2.03783697564280e+011 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port2_port6_p7 	_net_10 	gnd_0 	POLE 	_net_30 	gnd_0 	7.48954384169973e+009 	5.87361507022750e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010

* PORT_3
vi_3	port_3	_net_11	0.00000000000000e+000
vb_3	_net_14	_net_15	0.00000000000000e+000
R_Z0_3 	_net_11 	_net_12 	5.00000000000000e+001	NOISE=0
H_b_3	_net_12	gnd_0	vb_3	1.41421356237310e+001
E_v_3	_net_13	gnd_0	port_3	gnd_0	7.07106781186548e-002
H_i_3	_net_14	_net_13	vi_3	3.53553390593274e+000


G_POLE_port3_port1_p1 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	-3.65334497161625e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port3_port1_p2 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0  	3.72090655250536e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port3_port1_p3 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	-8.15745392526853e+008 	1.96340124318664e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port3_port1_p5 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	-4.01595725118987e+009 	-5.04466643655448e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port3_port1_p7 	_net_15 	gnd_0 	POLE 	_net_5 	gnd_0 	3.62923575837272e+009 	2.16260786971802e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port3_port2_p1 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	3.30221042406057e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port3_port2_p2 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0  	-1.51357824300096e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port3_port2_p3 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	-3.83896395732270e+008 	3.19628057927558e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port3_port2_p5 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	-7.96718679484474e+009 	5.50498003374687e+008 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port3_port2_p7 	_net_15 	gnd_0 	POLE 	_net_10 	gnd_0 	8.21479656290914e+009 	6.50142918198976e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port3_port3_p1 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.07490152233447e+008 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port3_port3_p2 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0  	1.83669540505128e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port3_port3_p3 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	-9.51007569487302e+008 	-1.60822251536047e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port3_port3_p5 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	-1.57111706981151e+010 	1.08537886151986e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port3_port3_p7 	_net_15 	gnd_0 	POLE 	_net_15 	gnd_0 	4.83052643091845e+009 	2.62351380093657e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port3_port4_p1 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	1.05576178818104e+008 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port3_port4_p2 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0  	-6.18756722891636e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port3_port4_p3 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	1.62842760492274e+010 	3.83913919322901e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port3_port4_p5 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	-8.54746244253431e+009 	-3.56176341321663e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port3_port4_p7 	_net_15 	gnd_0 	POLE 	_net_20 	gnd_0 	7.58072758870636e+009 	-3.11014808631771e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port3_port5_p1 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	-3.66924547035909e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port3_port5_p2 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0  	3.76495230947081e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port3_port5_p3 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.11300905300611e+009 	1.49824663942163e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port3_port5_p5 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	-4.23691059692524e+009 	-4.88989874983640e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port3_port5_p7 	_net_15 	gnd_0 	POLE 	_net_25 	gnd_0 	3.69792580308410e+009 	2.83019681679796e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port3_port6_p1 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	3.29613200742172e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port3_port6_p2 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.05899174200516e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port3_port6_p3 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	-6.41066168580740e+008 	2.00553845263024e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port3_port6_p5 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	-8.18783586600634e+009 	1.06169960223263e+008 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port3_port6_p7 	_net_15 	gnd_0 	POLE 	_net_30 	gnd_0 	8.25421907909966e+009 	6.74968962410325e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010

* PORT_4
vi_4	port_4	_net_16	0.00000000000000e+000
vb_4	_net_19	_net_20	0.00000000000000e+000
R_Z0_4 	_net_16 	_net_17 	5.00000000000000e+001	NOISE=0
H_b_4	_net_17	gnd_0	vb_4	1.41421356237310e+001
E_v_4	_net_18	gnd_0	port_4	gnd_0	7.07106781186548e-002
H_i_4	_net_19	_net_18	vi_4	3.53553390593274e+000


G_POLE_port4_port1_p1 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	3.32048496878048e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port4_port1_p2 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0  	-1.35988352969782e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port4_port1_p3 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	-3.29885451651886e+008 	3.69688277466882e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port4_port1_p5 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	-8.09091751240442e+009 	1.27427420869376e+009 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port4_port1_p7 	_net_20 	gnd_0 	POLE 	_net_5 	gnd_0 	8.14616163766072e+009 	6.65606949405473e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port4_port2_p1 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	-3.65578509876181e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port4_port2_p2 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0  	3.76406180657276e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port4_port2_p3 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.08800100515845e+009 	1.52634465650035e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port4_port2_p5 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	-4.25729105076331e+009 	-4.79159323433055e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port4_port2_p7 	_net_20 	gnd_0 	POLE 	_net_10 	gnd_0 	3.71033331149815e+009 	2.94237264253304e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port4_port3_p1 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	1.05576178818104e+008 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port4_port3_p2 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0  	-6.18756722891636e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port4_port3_p3 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	1.62842760492274e+010 	3.83913919322901e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port4_port3_p5 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	-8.54746244253431e+009 	-3.56176341321663e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port4_port3_p7 	_net_20 	gnd_0 	POLE 	_net_15 	gnd_0 	7.58072758870636e+009 	-3.11014808631771e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port4_port4_p1 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.07875754017829e+008 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port4_port4_p2 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0  	1.83257713529609e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port4_port4_p3 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.07080891987065e+009 	-1.40280567433601e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port4_port4_p5 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.58230681109063e+010 	1.00909929973939e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port4_port4_p7 	_net_20 	gnd_0 	POLE 	_net_20 	gnd_0 	4.66327787265166e+009 	2.69424343307097e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port4_port5_p1 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	3.28605366098291e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port4_port5_p2 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.09999298221112e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port4_port5_p3 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	-6.35140811098411e+008 	2.01822454189961e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port4_port5_p5 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	-8.13443455008975e+009 	1.99059584593010e+007 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port4_port5_p7 	_net_20 	gnd_0 	POLE 	_net_25 	gnd_0 	8.24178155224733e+009 	6.71128869279512e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port4_port6_p1 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	-3.69410008397164e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port4_port6_p2 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0  	3.79382558333373e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port4_port6_p3 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.38119636093789e+009 	1.24552077986315e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port4_port6_p5 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	-4.34535616618312e+009 	-4.85518619350632e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port4_port6_p7 	_net_20 	gnd_0 	POLE 	_net_30 	gnd_0 	3.75874348552333e+009 	3.38238198677969e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010

* PORT_5
vi_5	port_5	_net_21	0.00000000000000e+000
vb_5	_net_24	_net_25	0.00000000000000e+000
R_Z0_5 	_net_21 	_net_22 	5.00000000000000e+001	NOISE=0
H_b_5	_net_22	gnd_0	vb_5	1.41421356237310e+001
E_v_5	_net_23	gnd_0	port_5	gnd_0	7.07106781186548e-002
H_i_5	_net_24	_net_23	vi_5	3.53553390593274e+000


G_POLE_port5_port1_p1 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	2.38180432316301e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port5_port1_p2 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0  	2.39295455907431e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port5_port1_p3 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.05209892494071e+010 	2.57606540413510e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port5_port1_p5 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.12431904104578e+009 	-2.11874964036513e+011 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port5_port1_p7 	_net_25 	gnd_0 	POLE 	_net_5 	gnd_0 	7.55015440369252e+009 	5.56028200209978e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port5_port2_p1 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	-2.17049499682876e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port5_port2_p2 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0  	1.32455533654710e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port5_port2_p3 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-9.24479371195703e+009 	2.81748019695366e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port5_port2_p5 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.64409687181222e+009 	-8.61126622278852e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port5_port2_p7 	_net_25 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.16774917735257e+009 	-5.25465779412074e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port5_port3_p1 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	-3.66924547035909e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port5_port3_p2 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0  	3.76495230947081e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port5_port3_p3 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	-1.11300905300611e+009 	1.49824663942163e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port5_port3_p5 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	-4.23691059692524e+009 	-4.88989874983640e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port5_port3_p7 	_net_25 	gnd_0 	POLE 	_net_15 	gnd_0 	3.69792580308410e+009 	2.83019681679796e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port5_port4_p1 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	3.28605366098291e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port5_port4_p2 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0  	-1.09999298221112e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port5_port4_p3 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	-6.35140811098411e+008 	2.01822454189961e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port5_port4_p5 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	-8.13443455008975e+009 	1.99059584593010e+007 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port5_port4_p7 	_net_25 	gnd_0 	POLE 	_net_20 	gnd_0 	8.24178155224733e+009 	6.71128869279512e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port5_port5_p1 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	-8.54799855104162e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port5_port5_p2 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0  	6.76409391332339e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port5_port5_p3 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	7.56846791938578e+009 	4.45474853762058e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port5_port5_p5 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	-1.25051101071264e+010 	2.97346994131071e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port5_port5_p7 	_net_25 	gnd_0 	POLE 	_net_25 	gnd_0 	1.26241174461821e+009 	5.73333119580815e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port5_port6_p1 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	8.09462230414399e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port5_port6_p2 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0  	-1.14829434639448e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port5_port6_p3 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	2.22976495673276e+010 	3.33092960434431e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port5_port6_p5 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	-6.42438145700000e+009 	-2.87158598737472e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port5_port6_p7 	_net_25 	gnd_0 	POLE 	_net_30 	gnd_0 	4.81530185208258e+009 	-5.66056818725140e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010

* PORT_6
vi_6	port_6	_net_26	0.00000000000000e+000
vb_6	_net_29	_net_30	0.00000000000000e+000
R_Z0_6 	_net_26 	_net_27 	5.00000000000000e+001	NOISE=0
H_b_6	_net_27	gnd_0	vb_6	1.41421356237310e+001
E_v_6	_net_28	gnd_0	port_6	gnd_0	7.07106781186548e-002
H_i_6	_net_29	_net_28	vi_6	3.53553390593274e+000


G_POLE_port6_port1_p1 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	-2.14994539100996e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port6_port1_p2 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0  	1.34173277083232e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port6_port1_p3 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-9.22512997184087e+009 	2.82385839737405e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port6_port1_p5 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-2.78597977624556e+009 	-7.99222224234456e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port6_port1_p7 	_net_30 	gnd_0 	POLE 	_net_5 	gnd_0 	-1.21459579971251e+009 	-5.14290952085335e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port6_port2_p1 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	2.37875391275076e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port6_port2_p2 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0  	2.43560461434402e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port6_port2_p3 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	-1.08290404440687e+010 	2.55973078442315e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port6_port2_p5 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	-2.23526944528328e+009 	-2.03783697564280e+011 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port6_port2_p7 	_net_30 	gnd_0 	POLE 	_net_10 	gnd_0 	7.48954384169973e+009 	5.87361507022750e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port6_port3_p1 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	3.29613200742172e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port6_port3_p2 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0  	-1.05899174200516e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port6_port3_p3 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	-6.41066168580740e+008 	2.00553845263024e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port6_port3_p5 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	-8.18783586600634e+009 	1.06169960223263e+008 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port6_port3_p7 	_net_30 	gnd_0 	POLE 	_net_15 	gnd_0 	8.25421907909966e+009 	6.74968962410325e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port6_port4_p1 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	-3.69410008397164e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port6_port4_p2 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0  	3.79382558333373e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port6_port4_p3 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	-1.38119636093789e+009 	1.24552077986315e+011 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port6_port4_p5 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	-4.34535616618312e+009 	-4.85518619350632e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port6_port4_p7 	_net_30 	gnd_0 	POLE 	_net_20 	gnd_0 	3.75874348552333e+009 	3.38238198677969e+010 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port6_port5_p1 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	8.09462230414399e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port6_port5_p2 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0  	-1.14829434639448e+011 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port6_port5_p3 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	2.22976495673276e+010 	3.33092960434431e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port6_port5_p5 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	-6.42438145700000e+009 	-2.87158598737472e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port6_port5_p7 	_net_30 	gnd_0 	POLE 	_net_25 	gnd_0 	4.81530185208258e+009 	-5.66056818725140e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010
G_POLE_port6_port6_p1 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	-8.61082622569503e+007 / 1.0 	2.62516752593648e+009 , 0.0
G_POLE_port6_port6_p2 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0  	6.18768687660531e+010 / 1.0 	2.03878249406386e+012 , 0.0
G_POLE_port6_port6_p3 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	7.60545962027044e+009 	4.44533935560639e+010 , 0.0 / 1.0 	2.67197847788053e+010 , -8.26149049944623e+008
G_POLE_port6_port6_p5 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	-1.23631536008779e+010 	2.88726531389123e+010 , 0.0 / 1.0 	2.78552495029716e+010 , -5.26766780745907e+009
G_POLE_port6_port6_p7 	_net_30 	gnd_0 	POLE 	_net_30 	gnd_0 	1.14793651972439e+009 	5.97930653461207e+011 , 0.0 / 1.0 	3.01886130189647e+010 , -1.13594262644002e+010


.ENDS  bbspice_subckt
***************************************


***************************************
* S-based subckt

 
*bbspice subcircuit with external port numbers.

*.SUBCKT bbspice_Case4_10mm		1 	2 	3 	4 	5 	6 	0 

*x_ 	1 	2 	3 	4 	5 	6 	0 	bbspice_Case4_10mm_subckt

*.ENDS  bbspice_Case4_10mm
***************************************
*.ENDL
